`ifndef dut_interface_burst_config_v1_0_tb_include_vh_
`define dut_interface_burst_config_v1_0_tb_include_vh_

//Configuration current bd names
`define BD_INST_NAME dut_interface_burst_config_v1_0_bfm_1_i
`define BD_WRAPPER dut_interface_burst_config_v1_0_bfm_1_wrapper

//Configuration address parameters
`define S00_AXI_SLAVE_ADDRESS 32'h76000000
`define S01_AXI_SLAVE_ADDRESS 32'h44A00000
`endif
